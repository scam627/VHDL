----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:43:54 10/21/2017 
-- Design Name: 
-- Module Name:    SEU_IMM_MODULE - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SEU_IMM_MODULE is
    Port ( IMM : in  STD_LOGIC_VECTOR (12 downto 0);
           SIMM : out  STD_LOGIC_VECTOR (31 downto 0));
end SEU_IMM_MODULE;

architecture Behavioral of SEU_IMM_MODULE is

begin
	PROCESS(IMM)
	BEGIN
		CASE IMM(12) IS
			WHEN	'1' => SIMM <= STD_LOGIC_VECTOR("11111111111111111110000000000000"+IMM); 
			WHEN	OTHERS => SIMM <= STD_LOGIC_VECTOR("00000000000000000000000000000000"+IMM); 
		END CASE;
	END PROCESS;
end Behavioral;

